jbonepv
