module PU;
  logic [31:0]v1[7:0];  //1-D packed & 1-D unpacked (memory)
    
    initial begin
      //Array Index 7 of unpacked
      v1[7] = 'h FF_FF_FF_FF;  //equivalent to v1[7][31:0]
      
     
      
      
      //Array Index 6 of unpacked; 31:0 of packed
      v1[6][20:0] = 'h 11_11_11_11; 
      $display(v1);
      
      //Array Index 5 of unpacked; 15:0 of packed
      v1[5][15:0] = 'h aa_aa; 


      //Array Index 4 of unpacked; 0th bit of packed
      v1[4][0] = 1;  
      $display(v1);for(int i=7;i>=0;i--)
        for(int j=31;j>=0;j--)
          $display("value of v1[%0d][%0d] = %0d",i,j,v1[i][j]);
    end  
  endmodule
/*

# KERNEL: '{4294967295, X, x, x, x, x, x, x}
# KERNEL: '{4294967295, X, X, X, x, x, x, x}
# KERNEL: value of v1[7][31] = 1
# KERNEL: value of v1[7][30] = 1
# KERNEL: value of v1[7][29] = 1
# KERNEL: value of v1[7][28] = 1
# KERNEL: value of v1[7][27] = 1
# KERNEL: value of v1[7][26] = 1
# KERNEL: value of v1[7][25] = 1
# KERNEL: value of v1[7][24] = 1
# KERNEL: value of v1[7][23] = 1
# KERNEL: value of v1[7][22] = 1
# KERNEL: value of v1[7][21] = 1
# KERNEL: value of v1[7][20] = 1
# KERNEL: value of v1[7][19] = 1
# KERNEL: value of v1[7][18] = 1
# KERNEL: value of v1[7][17] = 1
# KERNEL: value of v1[7][16] = 1
# KERNEL: value of v1[7][15] = 1
# KERNEL: value of v1[7][14] = 1
# KERNEL: value of v1[7][13] = 1
# KERNEL: value of v1[7][12] = 1
# KERNEL: value of v1[7][11] = 1
# KERNEL: value of v1[7][10] = 1
# KERNEL: value of v1[7][9] = 1
# KERNEL: value of v1[7][8] = 1
# KERNEL: value of v1[7][7] = 1
# KERNEL: value of v1[7][6] = 1
# KERNEL: value of v1[7][5] = 1
# KERNEL: value of v1[7][4] = 1
# KERNEL: value of v1[7][3] = 1
# KERNEL: value of v1[7][2] = 1
# KERNEL: value of v1[7][1] = 1
# KERNEL: value of v1[7][0] = 1
# KERNEL: value of v1[6][31] = x
# KERNEL: value of v1[6][30] = x
# KERNEL: value of v1[6][29] = x
# KERNEL: value of v1[6][28] = x
# KERNEL: value of v1[6][27] = x
# KERNEL: value of v1[6][26] = x
# KERNEL: value of v1[6][25] = x
# KERNEL: value of v1[6][24] = x
# KERNEL: value of v1[6][23] = x
# KERNEL: value of v1[6][22] = x
# KERNEL: value of v1[6][21] = x
# KERNEL: value of v1[6][20] = 1
# KERNEL: value of v1[6][19] = 0
# KERNEL: value of v1[6][18] = 0
# KERNEL: value of v1[6][17] = 0
# KERNEL: value of v1[6][16] = 1
# KERNEL: value of v1[6][15] = 0
# KERNEL: value of v1[6][14] = 0
# KERNEL: value of v1[6][13] = 0
# KERNEL: value of v1[6][12] = 1
# KERNEL: value of v1[6][11] = 0
# KERNEL: value of v1[6][10] = 0
# KERNEL: value of v1[6][9] = 0
# KERNEL: value of v1[6][8] = 1
# KERNEL: value of v1[6][7] = 0
# KERNEL: value of v1[6][6] = 0
# KERNEL: value of v1[6][5] = 0
# KERNEL: value of v1[6][4] = 1
# KERNEL: value of v1[6][3] = 0
# KERNEL: value of v1[6][2] = 0
# KERNEL: value of v1[6][1] = 0
# KERNEL: value of v1[6][0] = 1
# KERNEL: value of v1[5][31] = x
# KERNEL: value of v1[5][30] = x
# KERNEL: value of v1[5][29] = x
# KERNEL: value of v1[5][28] = x
# KERNEL: value of v1[5][27] = x
# KERNEL: value of v1[5][26] = x
# KERNEL: value of v1[5][25] = x
# KERNEL: value of v1[5][24] = x
# KERNEL: value of v1[5][23] = x
# KERNEL: value of v1[5][22] = x
# KERNEL: value of v1[5][21] = x
# KERNEL: value of v1[5][20] = x
# KERNEL: value of v1[5][19] = x
# KERNEL: value of v1[5][18] = x
# KERNEL: value of v1[5][17] = x
# KERNEL: value of v1[5][16] = x
# KERNEL: value of v1[5][15] = 1
# KERNEL: value of v1[5][14] = 0
# KERNEL: value of v1[5][13] = 1
# KERNEL: value of v1[5][12] = 0
# KERNEL: value of v1[5][11] = 1
# KERNEL: value of v1[5][10] = 0
# KERNEL: value of v1[5][9] = 1
# KERNEL: value of v1[5][8] = 0
# KERNEL: value of v1[5][7] = 1
# KERNEL: value of v1[5][6] = 0
# KERNEL: value of v1[5][5] = 1
# KERNEL: value of v1[5][4] = 0
# KERNEL: value of v1[5][3] = 1
# KERNEL: value of v1[5][2] = 0
# KERNEL: value of v1[5][1] = 1
# KERNEL: value of v1[5][0] = 0
# KERNEL: value of v1[4][31] = x
# KERNEL: value of v1[4][30] = x
# KERNEL: value of v1[4][29] = x
# KERNEL: value of v1[4][28] = x
# KERNEL: value of v1[4][27] = x
# KERNEL: value of v1[4][26] = x
# KERNEL: value of v1[4][25] = x
# KERNEL: value of v1[4][24] = x
# KERNEL: value of v1[4][23] = x
# KERNEL: value of v1[4][22] = x
# KERNEL: value of v1[4][21] = x
# KERNEL: value of v1[4][20] = x
# KERNEL: value of v1[4][19] = x
# KERNEL: value of v1[4][18] = x
# KERNEL: value of v1[4][17] = x
# KERNEL: value of v1[4][16] = x
# KERNEL: value of v1[4][15] = x
# KERNEL: value of v1[4][14] = x
# KERNEL: value of v1[4][13] = x
# KERNEL: value of v1[4][12] = x
# KERNEL: value of v1[4][11] = x
# KERNEL: value of v1[4][10] = x
# KERNEL: value of v1[4][9] = x
# KERNEL: value of v1[4][8] = x
# KERNEL: value of v1[4][7] = x
# KERNEL: value of v1[4][6] = x
# KERNEL: value of v1[4][5] = x
# KERNEL: value of v1[4][4] = x
# KERNEL: value of v1[4][3] = x
# KERNEL: value of v1[4][2] = x
# KERNEL: value of v1[4][1] = x
# KERNEL: value of v1[4][0] = 1
# KERNEL: value of v1[3][31] = x
# KERNEL: value of v1[3][30] = x
# KERNEL: value of v1[3][29] = x
# KERNEL: value of v1[3][28] = x
# KERNEL: value of v1[3][27] = x
# KERNEL: value of v1[3][26] = x
# KERNEL: value of v1[3][25] = x
# KERNEL: value of v1[3][24] = x
# KERNEL: value of v1[3][23] = x
# KERNEL: value of v1[3][22] = x
# KERNEL: value of v1[3][21] = x
# KERNEL: value of v1[3][20] = x
# KERNEL: value of v1[3][19] = x
# KERNEL: value of v1[3][18] = x
# KERNEL: value of v1[3][17] = x
# KERNEL: value of v1[3][16] = x
# KERNEL: value of v1[3][15] = x
# KERNEL: value of v1[3][14] = x
# KERNEL: value of v1[3][13] = x
# KERNEL: value of v1[3][12] = x
# KERNEL: value of v1[3][11] = x
# KERNEL: value of v1[3][10] = x
# KERNEL: value of v1[3][9] = x
# KERNEL: value of v1[3][8] = x
# KERNEL: value of v1[3][7] = x
# KERNEL: value of v1[3][6] = x
# KERNEL: value of v1[3][5] = x
# KERNEL: value of v1[3][4] = x
# KERNEL: value of v1[3][3] = x
# KERNEL: value of v1[3][2] = x
# KERNEL: value of v1[3][1] = x
# KERNEL: value of v1[3][0] = x
# KERNEL: value of v1[2][31] = x
# KERNEL: value of v1[2][30] = x
# KERNEL: value of v1[2][29] = x
# KERNEL: value of v1[2][28] = x
# KERNEL: value of v1[2][27] = x
# KERNEL: value of v1[2][26] = x
# KERNEL: value of v1[2][25] = x
# KERNEL: value of v1[2][24] = x
# KERNEL: value of v1[2][23] = x
# KERNEL: value of v1[2][22] = x
# KERNEL: value of v1[2][21] = x
# KERNEL: value of v1[2][20] = x
# KERNEL: value of v1[2][19] = x
# KERNEL: value of v1[2][18] = x
# KERNEL: value of v1[2][17] = x
# KERNEL: value of v1[2][16] = x
# KERNEL: value of v1[2][15] = x
# KERNEL: value of v1[2][14] = x
# KERNEL: value of v1[2][13] = x
# KERNEL: value of v1[2][12] = x
# KERNEL: value of v1[2][11] = x
# KERNEL: value of v1[2][10] = x
# KERNEL: value of v1[2][9] = x
# KERNEL: value of v1[2][8] = x
# KERNEL: value of v1[2][7] = x
# KERNEL: value of v1[2][6] = x
# KERNEL: value of v1[2][5] = x
# KERNEL: value of v1[2][4] = x
# KERNEL: value of v1[2][3] = x
# KERNEL: value of v1[2][2] = x
# KERNEL: value of v1[2][1] = x
# KERNEL: value of v1[2][0] = x
# KERNEL: value of v1[1][31] = x
# KERNEL: value of v1[1][30] = x
# KERNEL: value of v1[1][29] = x
# KERNEL: value of v1[1][28] = x
# KERNEL: value of v1[1][27] = x
# KERNEL: value of v1[1][26] = x
# KERNEL: value of v1[1][25] = x
# KERNEL: value of v1[1][24] = x
# KERNEL: value of v1[1][23] = x
# KERNEL: value of v1[1][22] = x
# KERNEL: value of v1[1][21] = x
# KERNEL: value of v1[1][20] = x
# KERNEL: value of v1[1][19] = x
# KERNEL: value of v1[1][18] = x
# KERNEL: value of v1[1][17] = x
# KERNEL: value of v1[1][16] = x
# KERNEL: value of v1[1][15] = x
# KERNEL: value of v1[1][14] = x
# KERNEL: value of v1[1][13] = x
# KERNEL: value of v1[1][12] = x
# KERNEL: value of v1[1][11] = x
# KERNEL: value of v1[1][10] = x
# KERNEL: value of v1[1][9] = x
# KERNEL: value of v1[1][8] = x
# KERNEL: value of v1[1][7] = x
# KERNEL: value of v1[1][6] = x
# KERNEL: value of v1[1][5] = x
# KERNEL: value of v1[1][4] = x
# KERNEL: value of v1[1][3] = x
# KERNEL: value of v1[1][2] = x
# KERNEL: value of v1[1][1] = x
# KERNEL: value of v1[1][0] = x
# KERNEL: value of v1[0][31] = x
# KERNEL: value of v1[0][30] = x
# KERNEL: value of v1[0][29] = x
# KERNEL: value of v1[0][28] = x
# KERNEL: value of v1[0][27] = x
# KERNEL: value of v1[0][26] = x
# KERNEL: value of v1[0][25] = x
# KERNEL: value of v1[0][24] = x
# KERNEL: value of v1[0][23] = x
# KERNEL: value of v1[0][22] = x
# KERNEL: value of v1[0][21] = x
# KERNEL: value of v1[0][20] = x
# KERNEL: value of v1[0][19] = x
# KERNEL: value of v1[0][18] = x
# KERNEL: value of v1[0][17] = x
# KERNEL: value of v1[0][16] = x
# KERNEL: value of v1[0][15] = x
# KERNEL: value of v1[0][14] = x
# KERNEL: value of v1[0][13] = x
# KERNEL: value of v1[0][12] = x
# KERNEL: value of v1[0][11] = x
# KERNEL: value of v1[0][10] = x
# KERNEL: value of v1[0][9] = x
# KERNEL: value of v1[0][8] = x
# KERNEL: value of v1[0][7] = x
# KERNEL: value of v1[0][6] = x
# KERNEL: value of v1[0][5] = x
# KERNEL: value of v1[0][4] = x
# KERNEL: value of v1[0][3] = x
# KERNEL: value of v1[0][2] = x
# KERNEL: value of v1[0][1] = x
# KERNEL: value of v1[0][0] = x
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
# KERNEL: '{4294967295, X, x, x, x, x, x, x}
# KERNEL: '{4294967295, X, X, X, x, x, x, x}
# KERNEL: value of v1[7][31] = 1
# KERNEL: value of v1[7][30] = 1
# KERNEL: value of v1[7][29] = 1
# KERNEL: value of v1[7][28] = 1
# KERNEL: value of v1[7][27] = 1
# KERNEL: value of v1[7][26] = 1
# KERNEL: value of v1[7][25] = 1
# KERNEL: value of v1[7][24] = 1
# KERNEL: value of v1[7][23] = 1
# KERNEL: value of v1[7][22] = 1
# KERNEL: value of v1[7][21] = 1
# KERNEL: value of v1[7][20] = 1
# KERNEL: value of v1[7][19] = 1
# KERNEL: value of v1[7][18] = 1
# KERNEL: value of v1[7][17] = 1
# KERNEL: value of v1[7][16] = 1
# KERNEL: value of v1[7][15] = 1
# KERNEL: value of v1[7][14] = 1
# KERNEL: value of v1[7][13] = 1
# KERNEL: value of v1[7][12] = 1
# KERNEL: value of v1[7][11] = 1
# KERNEL: value of v1[7][10] = 1
# KERNEL: value of v1[7][9] = 1
# KERNEL: value of v1[7][8] = 1
# KERNEL: value of v1[7][7] = 1
# KERNEL: value of v1[7][6] = 1
# KERNEL: value of v1[7][5] = 1
# KERNEL: value of v1[7][4] = 1
# KERNEL: value of v1[7][3] = 1
# KERNEL: value of v1[7][2] = 1
# KERNEL: value of v1[7][1] = 1
# KERNEL: value of v1[7][0] = 1
# KERNEL: value of v1[6][31] = x
# KERNEL: value of v1[6][30] = x
# KERNEL: value of v1[6][29] = x
# KERNEL: value of v1[6][28] = x
# KERNEL: value of v1[6][27] = x
# KERNEL: value of v1[6][26] = x
# KERNEL: value of v1[6][25] = x
# KERNEL: value of v1[6][24] = x
# KERNEL: value of v1[6][23] = x
# KERNEL: value of v1[6][22] = x
# KERNEL: value of v1[6][21] = x
# KERNEL: value of v1[6][20] = 1
# KERNEL: value of v1[6][19] = 0
# KERNEL: value of v1[6][18] = 0
# KERNEL: value of v1[6][17] = 0
# KERNEL: value of v1[6][16] = 1
# KERNEL: value of v1[6][15] = 0
# KERNEL: value of v1[6][14] = 0
# KERNEL: value of v1[6][13] = 0
# KERNEL: value of v1[6][12] = 1
# KERNEL: value of v1[6][11] = 0
# KERNEL: value of v1[6][10] = 0
# KERNEL: value of v1[6][9] = 0
# KERNEL: value of v1[6][8] = 1
# KERNEL: value of v1[6][7] = 0
# KERNEL: value of v1[6][6] = 0
# KERNEL: value of v1[6][5] = 0
# KERNEL: value of v1[6][4] = 1
# KERNEL: value of v1[6][3] = 0
# KERNEL: value of v1[6][2] = 0
# KERNEL: value of v1[6][1] = 0
# KERNEL: value of v1[6][0] = 1
# KERNEL: value of v1[5][31] = x
# KERNEL: value of v1[5][30] = x
# KERNEL: value of v1[5][29] = x
# KERNEL: value of v1[5][28] = x
# KERNEL: value of v1[5][27] = x
# KERNEL: value of v1[5][26] = x
# KERNEL: value of v1[5][25] = x
# KERNEL: value of v1[5][24] = x
# KERNEL: value of v1[5][23] = x
# KERNEL: value of v1[5][22] = x
# KERNEL: value of v1[5][21] = x
# KERNEL: value of v1[5][20] = x
# KERNEL: value of v1[5][19] = x
# KERNEL: value of v1[5][18] = x
# KERNEL: value of v1[5][17] = x
# KERNEL: value of v1[5][16] = x
# KERNEL: value of v1[5][15] = 1
# KERNEL: value of v1[5][14] = 0
# KERNEL: value of v1[5][13] = 1
# KERNEL: value of v1[5][12] = 0
# KERNEL: value of v1[5][11] = 1
# KERNEL: value of v1[5][10] = 0
# KERNEL: value of v1[5][9] = 1
# KERNEL: value of v1[5][8] = 0
# KERNEL: value of v1[5][7] = 1
# KERNEL: value of v1[5][6] = 0
# KERNEL: value of v1[5][5] = 1
# KERNEL: value of v1[5][4] = 0
# KERNEL: value of v1[5][3] = 1
# KERNEL: value of v1[5][2] = 0
# KERNEL: value of v1[5][1] = 1
# KERNEL: value of v1[5][0] = 0
# KERNEL: value of v1[4][31] = x
# KERNEL: value of v1[4][30] = x
# KERNEL: value of v1[4][29] = x
# KERNEL: value of v1[4][28] = x
# KERNEL: value of v1[4][27] = x
# KERNEL: value of v1[4][26] = x
# KERNEL: value of v1[4][25] = x
# KERNEL: value of v1[4][24] = x
# KERNEL: value of v1[4][23] = x
# KERNEL: value of v1[4][22] = x
# KERNEL: value of v1[4][21] = x
# KERNEL: value of v1[4][20] = x
# KERNEL: value of v1[4][19] = x
# KERNEL: value of v1[4][18] = x
# KERNEL: value of v1[4][17] = x
# KERNEL: value of v1[4][16] = x
# KERNEL: value of v1[4][15] = x
# KERNEL: value of v1[4][14] = x
# KERNEL: value of v1[4][13] = x
# KERNEL: value of v1[4][12] = x
# KERNEL: value of v1[4][11] = x
# KERNEL: value of v1[4][10] = x
# KERNEL: value of v1[4][9] = x
# KERNEL: value of v1[4][8] = x
# KERNEL: value of v1[4][7] = x
# KERNEL: value of v1[4][6] = x
# KERNEL: value of v1[4][5] = x
# KERNEL: value of v1[4][4] = x
# KERNEL: value of v1[4][3] = x
# KERNEL: value of v1[4][2] = x
# KERNEL: value of v1[4][1] = x
# KERNEL: value of v1[4][0] = 1
# KERNEL: value of v1[3][31] = x
# KERNEL: value of v1[3][30] = x
# KERNEL: value of v1[3][29] = x
# KERNEL: value of v1[3][28] = x
# KERNEL: value of v1[3][27] = x
# KERNEL: value of v1[3][26] = x
# KERNEL: value of v1[3][25] = x
# KERNEL: value of v1[3][24] = x
# KERNEL: value of v1[3][23] = x
# KERNEL: value of v1[3][22] = x
# KERNEL: value of v1[3][21] = x
# KERNEL: value of v1[3][20] = x
# KERNEL: value of v1[3][19] = x
# KERNEL: value of v1[3][18] = x
# KERNEL: value of v1[3][17] = x
# KERNEL: value of v1[3][16] = x
# KERNEL: value of v1[3][15] = x
# KERNEL: value of v1[3][14] = x
# KERNEL: value of v1[3][13] = x
# KERNEL: value of v1[3][12] = x
# KERNEL: value of v1[3][11] = x
# KERNEL: value of v1[3][10] = x
# KERNEL: value of v1[3][9] = x
# KERNEL: value of v1[3][8] = x
# KERNEL: value of v1[3][7] = x
# KERNEL: value of v1[3][6] = x
# KERNEL: value of v1[3][5] = x
# KERNEL: value of v1[3][4] = x
# KERNEL: value of v1[3][3] = x
# KERNEL: value of v1[3][2] = x
# KERNEL: value of v1[3][1] = x
# KERNEL: value of v1[3][0] = x
# KERNEL: value of v1[2][31] = x
# KERNEL: value of v1[2][30] = x
# KERNEL: value of v1[2][29] = x
# KERNEL: value of v1[2][28] = x
# KERNEL: value of v1[2][27] = x
# KERNEL: value of v1[2][26] = x
# KERNEL: value of v1[2][25] = x
# KERNEL: value of v1[2][24] = x
# KERNEL: value of v1[2][23] = x
# KERNEL: value of v1[2][22] = x
# KERNEL: value of v1[2][21] = x
# KERNEL: value of v1[2][20] = x
# KERNEL: value of v1[2][19] = x
# KERNEL: value of v1[2][18] = x
# KERNEL: value of v1[2][17] = x
# KERNEL: value of v1[2][16] = x
# KERNEL: value of v1[2][15] = x
# KERNEL: value of v1[2][14] = x
# KERNEL: value of v1[2][13] = x
# KERNEL: value of v1[2][12] = x
# KERNEL: value of v1[2][11] = x
# KERNEL: value of v1[2][10] = x
# KERNEL: value of v1[2][9] = x
# KERNEL: value of v1[2][8] = x
# KERNEL: value of v1[2][7] = x
# KERNEL: value of v1[2][6] = x
# KERNEL: value of v1[2][5] = x
# KERNEL: value of v1[2][4] = x
# KERNEL: value of v1[2][3] = x
# KERNEL: value of v1[2][2] = x
# KERNEL: value of v1[2][1] = x
# KERNEL: value of v1[2][0] = x
# KERNEL: value of v1[1][31] = x
# KERNEL: value of v1[1][30] = x
# KERNEL: value of v1[1][29] = x
# KERNEL: value of v1[1][28] = x
# KERNEL: value of v1[1][27] = x
# KERNEL: value of v1[1][26] = x
# KERNEL: value of v1[1][25] = x
# KERNEL: value of v1[1][24] = x
# KERNEL: value of v1[1][23] = x
# KERNEL: value of v1[1][22] = x
# KERNEL: value of v1[1][21] = x
# KERNEL: value of v1[1][20] = x
# KERNEL: value of v1[1][19] = x
# KERNEL: value of v1[1][18] = x
# KERNEL: value of v1[1][17] = x
# KERNEL: value of v1[1][16] = x
# KERNEL: value of v1[1][15] = x
# KERNEL: value of v1[1][14] = x
# KERNEL: value of v1[1][13] = x
# KERNEL: value of v1[1][12] = x
# KERNEL: value of v1[1][11] = x
# KERNEL: value of v1[1][10] = x
# KERNEL: value of v1[1][9] = x
# KERNEL: value of v1[1][8] = x
# KERNEL: value of v1[1][7] = x
# KERNEL: value of v1[1][6] = x
# KERNEL: value of v1[1][5] = x
# KERNEL: value of v1[1][4] = x
# KERNEL: value of v1[1][3] = x
# KERNEL: value of v1[1][2] = x
# KERNEL: value of v1[1][1] = x
# KERNEL: value of v1[1][0] = x
# KERNEL: value of v1[0][31] = x
# KERNEL: value of v1[0][30] = x
# KERNEL: value of v1[0][29] = x
# KERNEL: value of v1[0][28] = x
# KERNEL: value of v1[0][27] = x
# KERNEL: value of v1[0][26] = x
# KERNEL: value of v1[0][25] = x
# KERNEL: value of v1[0][24] = x
# KERNEL: value of v1[0][23] = x
# KERNEL: value of v1[0][22] = x
# KERNEL: value of v1[0][21] = x
# KERNEL: value of v1[0][20] = x
# KERNEL: value of v1[0][19] = x
# KERNEL: value of v1[0][18] = x
# KERNEL: value of v1[0][17] = x
# KERNEL: value of v1[0][16] = x
# KERNEL: value of v1[0][15] = x
# KERNEL: value of v1[0][14] = x
# KERNEL: value of v1[0][13] = x
# KERNEL: value of v1[0][12] = x
# KERNEL: value of v1[0][11] = x
# KERNEL: value of v1[0][10] = x
# KERNEL: value of v1[0][9] = x
# KERNEL: value of v1[0][8] = x
# KERNEL: value of v1[0][7] = x
# KERNEL: value of v1[0][6] = x
# KERNEL: value of v1[0][5] = x
# KERNEL: value of v1[0][4] = x
# KERNEL: value of v1[0][3] = x
# KERNEL: value of v1[0][2] = x
# KERNEL: value of v1[0][1] = x
# KERNEL: value of v1[0][0] = x
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.

*/
