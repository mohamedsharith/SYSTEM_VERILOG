

`include "apb_2_i2c_defines.sv"
`include "apb_transaction.sv"
`include "apb_generator.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"


`include "i2c_transaction.sv"
`include "i2c_monitor.sv"
`include "apb_2_i2c_sb.sv"
`include "apb_2_i2c_env.sv"
`include "apb_2_i2c_test.sv"


