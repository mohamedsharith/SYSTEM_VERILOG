interface alu_int;  //don't use simply alu because we used that name in design so give a different name [error_spotted]
  logic a;
  logic b;
  logic alu_sel;
//   logic alu_expected;
  logic alu_out;
endinterface